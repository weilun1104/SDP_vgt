** Generated for: hspiceD
** Generated on: Mar 16 04:20:31 2024
** Design library name: ZYX_try
** Design cell name: bandgap_tb
** Design view name: schematic
.PARAM l1=0.6571um l2=2.7176um l3=5.9792um l4=2.0614um l5=0.5789um l6=4.1753um l7=1.4173um l8=2.6101um l9=1.8169um r1=3182944.0 r2=314825.8125 w1=14.9972um w2=49.6622um w3=84.1155um w4=20.5458um w5=2.5935um w6=14.9193um w7=40.8406um w8=20.1064um w9=38.3066um 



.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    HIER_DELIM=0

.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" BJT_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" DIO_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" RES_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" MIM_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" VAR_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" RES_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" MIM_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" VAR_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" IND_RF_PSUB_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" IND_RF_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 3TDIFF_PSUB_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 3TDIFF_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 2TDIFF_PSUB_TT
.LIB "C:\DAC\vanilla_bo_in_highdim-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 2TDIFF_TT

** Library name: ZYX_try
** Cell name: bandgap_1.8_v2
** View name: schematic
.subckt _sub3 gnd ib_ota vdd vref bias1 bias2
r7 _net0 net2 {r1}
r5 _net1 net1 {r1}
r4 net0136 _net1 {r2}
r0 net049 vref {r1}
q5 gnd gnd net049 pnp33a4 m=1
q4 gnd gnd _net0 pnp33a4 m=1
q3 gnd gnd net0136 pnp33a4 m=8
viprb0 sf_gate net021 DC=0
c8 sf_gate gnd mim w=25e-6 l=25e-6 m=8
m17 net030 bias1 net054 gnd n18 m=1 w=w4 l=l4 nf=6 ad='w4/6<419.5e-9?(int(3.0)*(176.4e-15+(w4/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w4/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w4/6))+(3.0-int(3.0)!=0?480e-9*(w4/6):0))/1' as='w4/6<419.5e-9?((((176.4e-15+(w4/6)*100e-9)+0*(w4/6<419.5e-9?420e-9:w4/6))+int(2.5)*(176.4e-15+(w4/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w4/6)*100e-9:0))/1:(((480e-9*(w4/6)+0*(w4/6<419.5e-9?420e-9:w4/6))+int(2.5)*(540e-9*(w4/6)))+(3.0-int(3.0)==0?480e-9*(w4/6):0))/1' pd='w4/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w4/6))+(3.0-int(3.0)!=0?960e-9+2*(w4/6):0))/1' ps='w4/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w4/6))+0)+int(2.5)*(1.08e-6+2*(w4/6)))+(3.0-int(3.0)==0?960e-9+2*(w4/6):0))/1' nrd='270e-9/((w4/6)*6)' nrs='270e-9/((w4/6)*6)' sa='w4/6<419.5e-9?520e-9:480e-9' sb='w4/6<419.5e-9?520e-9:480e-9' sd='w4/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
m14 net021 bias1 net055 gnd n18 m=1 w=w4 l=l4 nf=6 ad='w4/6<419.5e-9?(int(3.0)*(176.4e-15+(w4/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w4/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w4/6))+(3.0-int(3.0)!=0?480e-9*(w4/6):0))/1' as='w4/6<419.5e-9?((((176.4e-15+(w4/6)*100e-9)+0*(w4/6<419.5e-9?420e-9:w4/6))+int(2.5)*(176.4e-15+(w4/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w4/6)*100e-9:0))/1:(((480e-9*(w4/6)+0*(w4/6<419.5e-9?420e-9:w4/6))+int(2.5)*(540e-9*(w4/6)))+(3.0-int(3.0)==0?480e-9*(w4/6):0))/1' pd='w4/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w4/6))+(3.0-int(3.0)!=0?960e-9+2*(w4/6):0))/1' ps='w4/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w4/6))+0)+int(2.5)*(1.08e-6+2*(w4/6)))+(3.0-int(3.0)==0?960e-9+2*(w4/6):0))/1' nrd='270e-9/((w4/6)*6)' nrs='270e-9/((w4/6)*6)' sa='w4/6<419.5e-9?520e-9:480e-9' sb='w4/6<419.5e-9?520e-9:480e-9' sd='w4/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
m11 net055 _net0 net098 gnd n18 m=1 w=w5 l=l5 nf=4 ad='w5/4<419.5e-9?(int(2.0)*(176.4e-15+(w5/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w5/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w5/4))+(2.0-int(2.0)!=0?480e-9*(w5/4):0))/1' as='w5/4<419.5e-9?((((176.4e-15+(w5/4)*100e-9)+0*(w5/4<419.5e-9?420e-9:w5/4))+int(1.5)*(176.4e-15+(w5/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w5/4)*100e-9:0))/1:(((480e-9*(w5/4)+0*(w5/4<419.5e-9?420e-9:w5/4))+int(1.5)*(540e-9*(w5/4)))+(2.0-int(2.0)==0?480e-9*(w5/4):0))/1' pd='w5/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w5/4))+(2.0-int(2.0)!=0?960e-9+2*(w5/4):0))/1' ps='w5/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w5/4))+0)+int(1.5)*(1.08e-6+2*(w5/4)))+(2.0-int(2.0)==0?960e-9+2*(w5/4):0))/1' nrd='270e-9/((w5/4)*4)' nrs='270e-9/((w5/4)*4)' sa='w5/4<419.5e-9?520e-9:480e-9' sb='w5/4<419.5e-9?520e-9:480e-9' sd='w5/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
m10 net054 _net1 net098 gnd n18 m=1 w=w5 l=l5 nf=4 ad='w5/4<419.5e-9?(int(2.0)*(176.4e-15+(w5/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w5/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w5/4))+(2.0-int(2.0)!=0?480e-9*(w5/4):0))/1' as='w5/4<419.5e-9?((((176.4e-15+(w5/4)*100e-9)+0*(w5/4<419.5e-9?420e-9:w5/4))+int(1.5)*(176.4e-15+(w5/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w5/4)*100e-9:0))/1:(((480e-9*(w5/4)+0*(w5/4<419.5e-9?420e-9:w5/4))+int(1.5)*(540e-9*(w5/4)))+(2.0-int(2.0)==0?480e-9*(w5/4):0))/1' pd='w5/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w5/4))+(2.0-int(2.0)!=0?960e-9+2*(w5/4):0))/1' ps='w5/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w5/4))+0)+int(1.5)*(1.08e-6+2*(w5/4)))+(2.0-int(2.0)==0?960e-9+2*(w5/4):0))/1' nrd='270e-9/((w5/4)*4)' nrs='270e-9/((w5/4)*4)' sa='w5/4<419.5e-9?520e-9:480e-9' sb='w5/4<419.5e-9?520e-9:480e-9' sd='w5/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mnm4 bias1 bias1 bias2 gnd n18 m=1 w=w8 l=l8 nf=6 ad='w8/6<419.5e-9?(int(3.0)*(176.4e-15+(w8/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w8/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w8/6))+(3.0-int(3.0)!=0?480e-9*(w8/6):0))/1' as='w8/6<419.5e-9?((((176.4e-15+(w8/6)*100e-9)+0*(w8/6<419.5e-9?420e-9:w8/6))+int(2.5)*(176.4e-15+(w8/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w8/6)*100e-9:0))/1:(((480e-9*(w8/6)+0*(w8/6<419.5e-9?420e-9:w8/6))+int(2.5)*(540e-9*(w8/6)))+(3.0-int(3.0)==0?480e-9*(w8/6):0))/1' pd='w8/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w8/6))+(3.0-int(3.0)!=0?960e-9+2*(w8/6):0))/1' ps='w8/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w8/6))+0)+int(2.5)*(1.08e-6+2*(w8/6)))+(3.0-int(3.0)==0?960e-9+2*(w8/6):0))/1' nrd='270e-9/((w8/6)*6)' nrs='270e-9/((w8/6)*6)' sa='w8/6<419.5e-9?520e-9:480e-9' sb='w8/6<419.5e-9?520e-9:480e-9' sd='w8/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
m4 bias2 bias2 gnd gnd n18 m=1 w=w9 l=l9 nf=6 ad='w9/6<419.5e-9?(int(3.0)*(176.4e-15+(w9/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w9/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w9/6))+(3.0-int(3.0)!=0?480e-9*(w9/6):0))/1' as='w9/6<419.5e-9?((((176.4e-15+(w9/6)*100e-9)+0*(w9/6<419.5e-9?420e-9:w9/6))+int(2.5)*(176.4e-15+(w9/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w9/6)*100e-9:0))/1:(((480e-9*(w9/6)+0*(w9/6<419.5e-9?420e-9:w9/6))+int(2.5)*(540e-9*(w9/6)))+(3.0-int(3.0)==0?480e-9*(w9/6):0))/1' pd='w9/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w9/6))+(3.0-int(3.0)!=0?960e-9+2*(w9/6):0))/1' ps='w9/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w9/6))+0)+int(2.5)*(1.08e-6+2*(w9/6)))+(3.0-int(3.0)==0?960e-9+2*(w9/6):0))/1' nrd='270e-9/((w9/6)*6)' nrs='270e-9/((w9/6)*6)' sa='w9/6<419.5e-9?520e-9:480e-9' sb='w9/6<419.5e-9?520e-9:480e-9' sd='w9/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
m3 net098 bias2 gnd gnd n18 m=1 w=w6 l=l6 nf=6 ad='w6/6<419.5e-9?(int(3.0)*(176.4e-15+(w6/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w6/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w6/6))+(3.0-int(3.0)!=0?480e-9*(w6/6):0))/1' as='w6/6<419.5e-9?((((176.4e-15+(w6/6)*100e-9)+0*(w6/6<419.5e-9?420e-9:w6/6))+int(2.5)*(176.4e-15+(w6/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w6/6)*100e-9:0))/1:(((480e-9*(w6/6)+0*(w6/6<419.5e-9?420e-9:w6/6))+int(2.5)*(540e-9*(w6/6)))+(3.0-int(3.0)==0?480e-9*(w6/6):0))/1' pd='w6/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w6/6))+(3.0-int(3.0)!=0?960e-9+2*(w6/6):0))/1' ps='w6/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w6/6))+0)+int(2.5)*(1.08e-6+2*(w6/6)))+(3.0-int(3.0)==0?960e-9+2*(w6/6):0))/1' nrd='270e-9/((w6/6)*6)' nrs='270e-9/((w6/6)*6)' sa='w6/6<419.5e-9?520e-9:480e-9' sb='w6/6<419.5e-9?520e-9:480e-9' sd='w6/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm56 net6 net6 vdd vdd p18 m=1 w=30e-6 l=1e-6 nf=1 ad=14.4e-12 as=14.4e-12 pd=60.96e-6 ps=60.96e-6 nrd=9e-3 nrs=9e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mpm55 net3 net3 vdd vdd p18 m=1 w=30e-6 l=1e-6 nf=1 ad=14.4e-12 as=14.4e-12 pd=60.96e-6 ps=60.96e-6 nrd=9e-3 nrs=9e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mpm54 net4 net4 vdd vdd p18 m=1 w=30e-6 l=1e-6 nf=1 ad=14.4e-12 as=14.4e-12 pd=60.96e-6 ps=60.96e-6 nrd=9e-3 nrs=9e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mpm53 net5 net5 vdd vdd p18 m=1 w=30e-6 l=1e-6 nf=1 ad=14.4e-12 as=14.4e-12 pd=60.96e-6 ps=60.96e-6 nrd=9e-3 nrs=9e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mpm19 net1 sf_gate net5 net5 p18 m=1 w=w1 l=l1 nf=1 ad='w1/1<419.5e-9?(int(500e-3)*(176.4e-15+(w1/1)*200e-9)+(500e-3-int(500e-3)!=0?176.4e-15+(w1/1)*100e-9:0))/1:(int(500e-3)*(540e-9*(w1/1))+(500e-3-int(500e-3)!=0?480e-9*(w1/1):0))/1' as='w1/1<419.5e-9?((((176.4e-15+(w1/1)*100e-9)+0*(w1/1<419.5e-9?420e-9:w1/1))+int(0.0)*(176.4e-15+(w1/1)*200e-9))+(500e-3-int(500e-3)==0?176.4e-15+(w1/1)*100e-9:0))/1:(((480e-9*(w1/1)+0*(w1/1<419.5e-9?420e-9:w1/1))+int(0.0)*(540e-9*(w1/1)))+(500e-3-int(500e-3)==0?480e-9*(w1/1):0))/1' pd='w1/1<419.5e-9?(int(500e-3)*2.08e-6+(500e-3-int(500e-3)!=0?1.88e-6:0))/1:(int(500e-3)*(1.08e-6+2*(w1/1))+(500e-3-int(500e-3)!=0?960e-9+2*(w1/1):0))/1' ps='w1/1<419.5e-9?((1.88e-6+int(0.0)*2.08e-6)+(500e-3-int(500e-3)==0?1.88e-6:0))/1:((((960e-9+2*(w1/1))+0)+int(0.0)*(1.08e-6+2*(w1/1)))+(500e-3-int(500e-3)==0?960e-9+2*(w1/1):0))/1' nrd='270e-9/((w1/1)*1)' nrs='270e-9/((w1/1)*1)' sa='w1/1<419.5e-9?520e-9:480e-9' sb='w1/1<419.5e-9?520e-9:480e-9' sd=0 sca=0 scb=0 scc=0
mpm20 ib_ota sf_gate net6 net6 p18 m=1 w=w1 l=l1 nf=1 ad='w1/1<419.5e-9?(int(500e-3)*(176.4e-15+(w1/1)*200e-9)+(500e-3-int(500e-3)!=0?176.4e-15+(w1/1)*100e-9:0))/1:(int(500e-3)*(540e-9*(w1/1))+(500e-3-int(500e-3)!=0?480e-9*(w1/1):0))/1' as='w1/1<419.5e-9?((((176.4e-15+(w1/1)*100e-9)+0*(w1/1<419.5e-9?420e-9:w1/1))+int(0.0)*(176.4e-15+(w1/1)*200e-9))+(500e-3-int(500e-3)==0?176.4e-15+(w1/1)*100e-9:0))/1:(((480e-9*(w1/1)+0*(w1/1<419.5e-9?420e-9:w1/1))+int(0.0)*(540e-9*(w1/1)))+(500e-3-int(500e-3)==0?480e-9*(w1/1):0))/1' pd='w1/1<419.5e-9?(int(500e-3)*2.08e-6+(500e-3-int(500e-3)!=0?1.88e-6:0))/1:(int(500e-3)*(1.08e-6+2*(w1/1))+(500e-3-int(500e-3)!=0?960e-9+2*(w1/1):0))/1' ps='w1/1<419.5e-9?((1.88e-6+int(0.0)*2.08e-6)+(500e-3-int(500e-3)==0?1.88e-6:0))/1:((((960e-9+2*(w1/1))+0)+int(0.0)*(1.08e-6+2*(w1/1)))+(500e-3-int(500e-3)==0?960e-9+2*(w1/1):0))/1' nrd='270e-9/((w1/1)*1)' nrs='270e-9/((w1/1)*1)' sa='w1/1<419.5e-9?520e-9:480e-9' sb='w1/1<419.5e-9?520e-9:480e-9' sd=0 sca=0 scb=0 scc=0
m25 net021 net030 net020 net020 p18 m=1 w=w3 l=l3 nf=6 ad='w3/6<419.5e-9?(int(3.0)*(176.4e-15+(w3/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w3/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w3/6))+(3.0-int(3.0)!=0?480e-9*(w3/6):0))/1' as='w3/6<419.5e-9?((((176.4e-15+(w3/6)*100e-9)+0*(w3/6<419.5e-9?420e-9:w3/6))+int(2.5)*(176.4e-15+(w3/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w3/6)*100e-9:0))/1:(((480e-9*(w3/6)+0*(w3/6<419.5e-9?420e-9:w3/6))+int(2.5)*(540e-9*(w3/6)))+(3.0-int(3.0)==0?480e-9*(w3/6):0))/1' pd='w3/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w3/6))+(3.0-int(3.0)!=0?960e-9+2*(w3/6):0))/1' ps='w3/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w3/6))+0)+int(2.5)*(1.08e-6+2*(w3/6)))+(3.0-int(3.0)==0?960e-9+2*(w3/6):0))/1' nrd='270e-9/((w3/6)*6)' nrs='270e-9/((w3/6)*6)' sa='w3/6<419.5e-9?520e-9:480e-9' sb='w3/6<419.5e-9?520e-9:480e-9' sd='w3/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
m24 net030 net030 net025 net025 p18 m=1 w=w3 l=l3 nf=6 ad='w3/6<419.5e-9?(int(3.0)*(176.4e-15+(w3/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w3/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w3/6))+(3.0-int(3.0)!=0?480e-9*(w3/6):0))/1' as='w3/6<419.5e-9?((((176.4e-15+(w3/6)*100e-9)+0*(w3/6<419.5e-9?420e-9:w3/6))+int(2.5)*(176.4e-15+(w3/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w3/6)*100e-9:0))/1:(((480e-9*(w3/6)+0*(w3/6<419.5e-9?420e-9:w3/6))+int(2.5)*(540e-9*(w3/6)))+(3.0-int(3.0)==0?480e-9*(w3/6):0))/1' pd='w3/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w3/6))+(3.0-int(3.0)!=0?960e-9+2*(w3/6):0))/1' ps='w3/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w3/6))+0)+int(2.5)*(1.08e-6+2*(w3/6)))+(3.0-int(3.0)==0?960e-9+2*(w3/6):0))/1' nrd='270e-9/((w3/6)*6)' nrs='270e-9/((w3/6)*6)' sa='w3/6<419.5e-9?520e-9:480e-9' sb='w3/6<419.5e-9?520e-9:480e-9' sd='w3/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm24 net2 sf_gate net4 net4 p18 m=1 w=w1 l=l1 nf=1 ad='w1/1<419.5e-9?(int(500e-3)*(176.4e-15+(w1/1)*200e-9)+(500e-3-int(500e-3)!=0?176.4e-15+(w1/1)*100e-9:0))/1:(int(500e-3)*(540e-9*(w1/1))+(500e-3-int(500e-3)!=0?480e-9*(w1/1):0))/1' as='w1/1<419.5e-9?((((176.4e-15+(w1/1)*100e-9)+0*(w1/1<419.5e-9?420e-9:w1/1))+int(0.0)*(176.4e-15+(w1/1)*200e-9))+(500e-3-int(500e-3)==0?176.4e-15+(w1/1)*100e-9:0))/1:(((480e-9*(w1/1)+0*(w1/1<419.5e-9?420e-9:w1/1))+int(0.0)*(540e-9*(w1/1)))+(500e-3-int(500e-3)==0?480e-9*(w1/1):0))/1' pd='w1/1<419.5e-9?(int(500e-3)*2.08e-6+(500e-3-int(500e-3)!=0?1.88e-6:0))/1:(int(500e-3)*(1.08e-6+2*(w1/1))+(500e-3-int(500e-3)!=0?960e-9+2*(w1/1):0))/1' ps='w1/1<419.5e-9?((1.88e-6+int(0.0)*2.08e-6)+(500e-3-int(500e-3)==0?1.88e-6:0))/1:((((960e-9+2*(w1/1))+0)+int(0.0)*(1.08e-6+2*(w1/1)))+(500e-3-int(500e-3)==0?960e-9+2*(w1/1):0))/1' nrd='270e-9/((w1/1)*1)' nrs='270e-9/((w1/1)*1)' sa='w1/1<419.5e-9?520e-9:480e-9' sb='w1/1<419.5e-9?520e-9:480e-9' sd=0 sca=0 scb=0 scc=0
mpm31 net025 net025 vdd vdd p18 m=1 w=w2 l=l2 nf=6 ad='w2/6<419.5e-9?(int(3.0)*(176.4e-15+(w2/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w2/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w2/6))+(3.0-int(3.0)!=0?480e-9*(w2/6):0))/1' as='w2/6<419.5e-9?((((176.4e-15+(w2/6)*100e-9)+0*(w2/6<419.5e-9?420e-9:w2/6))+int(2.5)*(176.4e-15+(w2/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w2/6)*100e-9:0))/1:(((480e-9*(w2/6)+0*(w2/6<419.5e-9?420e-9:w2/6))+int(2.5)*(540e-9*(w2/6)))+(3.0-int(3.0)==0?480e-9*(w2/6):0))/1' pd='w2/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w2/6))+(3.0-int(3.0)!=0?960e-9+2*(w2/6):0))/1' ps='w2/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w2/6))+0)+int(2.5)*(1.08e-6+2*(w2/6)))+(3.0-int(3.0)==0?960e-9+2*(w2/6):0))/1' nrd='270e-9/((w2/6)*6)' nrs='270e-9/((w2/6)*6)' sa='w2/6<419.5e-9?520e-9:480e-9' sb='w2/6<419.5e-9?520e-9:480e-9' sd='w2/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm32 net020 net025 vdd vdd p18 m=1 w=w2 l=l2 nf=6 ad='w2/6<419.5e-9?(int(3.0)*(176.4e-15+(w2/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w2/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w2/6))+(3.0-int(3.0)!=0?480e-9*(w2/6):0))/1' as='w2/6<419.5e-9?((((176.4e-15+(w2/6)*100e-9)+0*(w2/6<419.5e-9?420e-9:w2/6))+int(2.5)*(176.4e-15+(w2/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w2/6)*100e-9:0))/1:(((480e-9*(w2/6)+0*(w2/6<419.5e-9?420e-9:w2/6))+int(2.5)*(540e-9*(w2/6)))+(3.0-int(3.0)==0?480e-9*(w2/6):0))/1' pd='w2/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w2/6))+(3.0-int(3.0)!=0?960e-9+2*(w2/6):0))/1' ps='w2/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w2/6))+0)+int(2.5)*(1.08e-6+2*(w2/6)))+(3.0-int(3.0)==0?960e-9+2*(w2/6):0))/1' nrd='270e-9/((w2/6)*6)' nrs='270e-9/((w2/6)*6)' sa='w2/6<419.5e-9?520e-9:480e-9' sb='w2/6<419.5e-9?520e-9:480e-9' sd='w2/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm21 vref sf_gate net3 net3 p18 m=1 w=w1 l=l1 nf=1 ad='w1/1<419.5e-9?(int(500e-3)*(176.4e-15+(w1/1)*200e-9)+(500e-3-int(500e-3)!=0?176.4e-15+(w1/1)*100e-9:0))/1:(int(500e-3)*(540e-9*(w1/1))+(500e-3-int(500e-3)!=0?480e-9*(w1/1):0))/1' as='w1/1<419.5e-9?((((176.4e-15+(w1/1)*100e-9)+0*(w1/1<419.5e-9?420e-9:w1/1))+int(0.0)*(176.4e-15+(w1/1)*200e-9))+(500e-3-int(500e-3)==0?176.4e-15+(w1/1)*100e-9:0))/1:(((480e-9*(w1/1)+0*(w1/1<419.5e-9?420e-9:w1/1))+int(0.0)*(540e-9*(w1/1)))+(500e-3-int(500e-3)==0?480e-9*(w1/1):0))/1' pd='w1/1<419.5e-9?(int(500e-3)*2.08e-6+(500e-3-int(500e-3)!=0?1.88e-6:0))/1:(int(500e-3)*(1.08e-6+2*(w1/1))+(500e-3-int(500e-3)!=0?960e-9+2*(w1/1):0))/1' ps='w1/1<419.5e-9?((1.88e-6+int(0.0)*2.08e-6)+(500e-3-int(500e-3)==0?1.88e-6:0))/1:((((960e-9+2*(w1/1))+0)+int(0.0)*(1.08e-6+2*(w1/1)))+(500e-3-int(500e-3)==0?960e-9+2*(w1/1):0))/1' nrd='270e-9/((w1/1)*1)' nrs='270e-9/((w1/1)*1)' sa='w1/1<419.5e-9?520e-9:480e-9' sb='w1/1<419.5e-9?520e-9:480e-9' sd=0 sca=0 scb=0 scc=0
mpm33 bias1 bias1 vdd vdd p18 m=1 w=w7 l=l7 nf=6 ad='w7/6<419.5e-9?(int(3.0)*(176.4e-15+(w7/6)*200e-9)+(3.0-int(3.0)!=0?176.4e-15+(w7/6)*100e-9:0))/1:(int(3.0)*(540e-9*(w7/6))+(3.0-int(3.0)!=0?480e-9*(w7/6):0))/1' as='w7/6<419.5e-9?((((176.4e-15+(w7/6)*100e-9)+0*(w7/6<419.5e-9?420e-9:w7/6))+int(2.5)*(176.4e-15+(w7/6)*200e-9))+(3.0-int(3.0)==0?176.4e-15+(w7/6)*100e-9:0))/1:(((480e-9*(w7/6)+0*(w7/6<419.5e-9?420e-9:w7/6))+int(2.5)*(540e-9*(w7/6)))+(3.0-int(3.0)==0?480e-9*(w7/6):0))/1' pd='w7/6<419.5e-9?(int(3.0)*2.08e-6+(3.0-int(3.0)!=0?1.88e-6:0))/1:(int(3.0)*(1.08e-6+2*(w7/6))+(3.0-int(3.0)!=0?960e-9+2*(w7/6):0))/1' ps='w7/6<419.5e-9?((1.88e-6+int(2.5)*2.08e-6)+(3.0-int(3.0)==0?1.88e-6:0))/1:((((960e-9+2*(w7/6))+0)+int(2.5)*(1.08e-6+2*(w7/6)))+(3.0-int(3.0)==0?960e-9+2*(w7/6):0))/1' nrd='270e-9/((w7/6)*6)' nrs='270e-9/((w7/6)*6)' sa='w7/6<419.5e-9?520e-9:480e-9' sb='w7/6<419.5e-9?520e-9:480e-9' sd='w7/6<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
.ends _sub3
** End of subcircuit definition.

** Library name: ZYX_try
** Cell name: bandgap_tb
** View name: schematic
xi17 0 net3 vdd vref net8 net9 _sub3
r2 net3 0 1e6
v0 vdd 0 DC=1.8 AC 1

.control
op
dc TEMP -40 125 1
ac dec 10 1 100000K
ac lin 1 1 2
.endc

.END
