** Generated for: hspiceD
** Generated on: Jan 26 20:27:58 2024
** Design library name: ZYX_try
** Design cell name: 5_T_OTA_tb
** Design view name: schematic
.PARAM l1=1.5611271890610412e-06 l2=4.934858792566221e-06 l3=6.884146555959352e-07 w1=0.00017482827972199695 w2=0.00011018140467152217 w3=4.9892637417140984e-05  



.AC DEC 10  

.DC    

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    HIER_DELIM=0
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" BJT_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" DIO_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" RES_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" MIM_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" VAR_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" RES_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" MIM_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" VAR_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" IND_RF_PSUB_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" IND_RF_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 3TDIFF_PSUB_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 3TDIFF_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 2TDIFF_PSUB_TT
.LIB "C:\Users\icelab01\Desktop\ZhuohuaLiu_2024_BYA_jiebang\BYA_jiebang\BYA_jiebang\Knowledge_unbinding\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 2TDIFF_TT

** Library name: ZYX_try
** Cell name: 5_T_OTA
** View name: schematic
.subckt ZYX_try_5_T_OTA_schematic gnd iss vn vout vp vss
mpm1 vss net2 vout vss p18 m=1 w=w2 l=l2 nf=4 ad='w2/4<419.5e-9?(int(2.0)*(176.4e-15+(w2/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w2/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w2/4))+(2.0-int(2.0)!=0?480e-9*(w2/4):0))/1' as='w2/4<419.5e-9?((((176.4e-15+(w2/4)*100e-9)+0*(w2/4<419.5e-9?420e-9:w2/4))+int(1.5)*(176.4e-15+(w2/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w2/4)*100e-9:0))/1:(((480e-9*(w2/4)+0*(w2/4<419.5e-9?420e-9:w2/4))+int(1.5)*(540e-9*(w2/4)))+(2.0-int(2.0)==0?480e-9*(w2/4):0))/1' pd='w2/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w2/4))+(2.0-int(2.0)!=0?960e-9+2*(w2/4):0))/1' ps='w2/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w2/4))+0)+int(1.5)*(1.08e-6+2*(w2/4)))+(2.0-int(2.0)==0?960e-9+2*(w2/4):0))/1' nrd='270e-9/((w2/4)*4)' nrs='270e-9/((w2/4)*4)' sa='w2/4<419.5e-9?520e-9:480e-9' sb='w2/4<419.5e-9?520e-9:480e-9' sd='w2/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm0 net2 net2 vss vss p18 m=1 w=w2 l=l2 nf=4 ad='w2/4<419.5e-9?(int(2.0)*(176.4e-15+(w2/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w2/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w2/4))+(2.0-int(2.0)!=0?480e-9*(w2/4):0))/1' as='w2/4<419.5e-9?((((176.4e-15+(w2/4)*100e-9)+0*(w2/4<419.5e-9?420e-9:w2/4))+int(1.5)*(176.4e-15+(w2/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w2/4)*100e-9:0))/1:(((480e-9*(w2/4)+0*(w2/4<419.5e-9?420e-9:w2/4))+int(1.5)*(540e-9*(w2/4)))+(2.0-int(2.0)==0?480e-9*(w2/4):0))/1' pd='w2/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w2/4))+(2.0-int(2.0)!=0?960e-9+2*(w2/4):0))/1' ps='w2/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w2/4))+0)+int(1.5)*(1.08e-6+2*(w2/4)))+(2.0-int(2.0)==0?960e-9+2*(w2/4):0))/1' nrd='270e-9/((w2/4)*4)' nrs='270e-9/((w2/4)*4)' sa='w2/4<419.5e-9?520e-9:480e-9' sb='w2/4<419.5e-9?520e-9:480e-9' sd='w2/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mnm7 iss iss gnd gnd n18 m=1 w=130e-6 l=1e-6 nf=4 ad=35.1e-12 as=48.75e-12 pd=132.16e-6 ps=198e-6 nrd=2.07692e-3 nrs=2.07692e-3 sa=480e-9 sb=480e-9 sd=540e-9 sca=0 scb=0 scc=0
mnm2 net1 iss gnd gnd n18 m=1 w=w3 l=l3 nf=4 ad='w3/4<419.5e-9?(int(2.0)*(176.4e-15+(w3/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w3/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w3/4))+(2.0-int(2.0)!=0?480e-9*(w3/4):0))/1' as='w3/4<419.5e-9?((((176.4e-15+(w3/4)*100e-9)+0*(w3/4<419.5e-9?420e-9:w3/4))+int(1.5)*(176.4e-15+(w3/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w3/4)*100e-9:0))/1:(((480e-9*(w3/4)+0*(w3/4<419.5e-9?420e-9:w3/4))+int(1.5)*(540e-9*(w3/4)))+(2.0-int(2.0)==0?480e-9*(w3/4):0))/1' pd='w3/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w3/4))+(2.0-int(2.0)!=0?960e-9+2*(w3/4):0))/1' ps='w3/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w3/4))+0)+int(1.5)*(1.08e-6+2*(w3/4)))+(2.0-int(2.0)==0?960e-9+2*(w3/4):0))/1' nrd='270e-9/((w3/4)*4)' nrs='270e-9/((w3/4)*4)' sa='w3/4<419.5e-9?520e-9:480e-9' sb='w3/4<419.5e-9?520e-9:480e-9' sd='w3/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mnm1 net1 vn vout gnd n18 m=1 w=w1 l=l1 nf=4 ad='w1/4<419.5e-9?(int(2.0)*(176.4e-15+(w1/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w1/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w1/4))+(2.0-int(2.0)!=0?480e-9*(w1/4):0))/1' as='w1/4<419.5e-9?((((176.4e-15+(w1/4)*100e-9)+0*(w1/4<419.5e-9?420e-9:w1/4))+int(1.5)*(176.4e-15+(w1/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w1/4)*100e-9:0))/1:(((480e-9*(w1/4)+0*(w1/4<419.5e-9?420e-9:w1/4))+int(1.5)*(540e-9*(w1/4)))+(2.0-int(2.0)==0?480e-9*(w1/4):0))/1' pd='w1/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w1/4))+(2.0-int(2.0)!=0?960e-9+2*(w1/4):0))/1' ps='w1/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w1/4))+0)+int(1.5)*(1.08e-6+2*(w1/4)))+(2.0-int(2.0)==0?960e-9+2*(w1/4):0))/1' nrd='270e-9/((w1/4)*4)' nrs='270e-9/((w1/4)*4)' sa='w1/4<419.5e-9?520e-9:480e-9' sb='w1/4<419.5e-9?520e-9:480e-9' sd='w1/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mnm0 net2 vp net1 gnd n18 m=1 w=w1 l=l1 nf=4 ad='w1/4<419.5e-9?(int(2.0)*(176.4e-15+(w1/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w1/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w1/4))+(2.0-int(2.0)!=0?480e-9*(w1/4):0))/1' as='w1/4<419.5e-9?((((176.4e-15+(w1/4)*100e-9)+0*(w1/4<419.5e-9?420e-9:w1/4))+int(1.5)*(176.4e-15+(w1/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w1/4)*100e-9:0))/1:(((480e-9*(w1/4)+0*(w1/4<419.5e-9?420e-9:w1/4))+int(1.5)*(540e-9*(w1/4)))+(2.0-int(2.0)==0?480e-9*(w1/4):0))/1' pd='w1/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w1/4))+(2.0-int(2.0)!=0?960e-9+2*(w1/4):0))/1' ps='w1/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w1/4))+0)+int(1.5)*(1.08e-6+2*(w1/4)))+(2.0-int(2.0)==0?960e-9+2*(w1/4):0))/1' nrd='270e-9/((w1/4)*4)' nrs='270e-9/((w1/4)*4)' sa='w1/4<419.5e-9?520e-9:480e-9' sb='w1/4<419.5e-9?520e-9:480e-9' sd='w1/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
.ends ZYX_try_5_T_OTA_schematic
** End of subcircuit definition.

** Library name: ZYX_try
** Cell name: 5_T_OTA_tb
** View name: schematic
xi3 0 iss net2 net3 net1 vss ZYX_try_5_T_OTA_schematic
v8 vss 0 DC=3.3 AC 0
v1 net1 0 DC=1.65 AC 0
v0 net2 net1 DC=0 AC 1 180
c0 net3 0 5e-12
i4 vss iss DC=1e-3

.control
op
AC DEC 10 0.01 100000K
settype decibel out
plot vdb(net3) xlimit 1 100000k ylabel 'small signal gain'
settype phase out
plot cph(net3) xlimit 1 100000k ylabel 'phase (in rad)'
let outd = 180/PI*cph(net3)
settype phase outd
plot outd xlimit 1 100000k ylabel 'phase'
.endc

.END
