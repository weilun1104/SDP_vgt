** Generated for: hspiceD
** Generated on: Mar  1 08:28:19 2024
** Design library name: ZYX_try
** Design cell name: tb_OTA_three
** Design view name: schematic
.GLOBAL vdd!
.PARAM c1=5.73pf c2=3.04pf l1=0.83u l2=0.47u l3=0.94u l4=1.94u l5=0.95u l6=0.61u l7=1.09u l8=1.14u w1=5.28u w2=2.57u w3=75.37u w4=35.04u w5=3.67u w6=5.22u w7=68.16u w8=124.36u



.PROBE DC
+    V(net1)
+    V(net2)
.PROBE AC
+    V(net1) VP(net1)
+    V(net2) VP(net2)
.AC DEC 10  

.DC    

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
+    HIER_DELIM=0
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" BJT_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" DIO_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" RES_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" MIM_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\ms018_enhanced_v1p11.lib" VAR_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" RES_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" MIM_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" VAR_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" IND_RF_PSUB_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" IND_RF_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 3TDIFF_PSUB_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 3TDIFF_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 2TDIFF_PSUB_TT
.LIB "C:\DAC\VGT-main\Simulation\Data\smic18\models\hspice\mse018_v1p11_rf.lib" 2TDIFF_TT

** Library name: yaoyuan
** Cell name: OTA_three
** View name: schematic
.subckt OTA_three _net1 _net0 vout
mnm6 bias1 bias1 0 0 n18 m=1 w=3e-6 l=1e-6 nf=1 ad=1.44e-12 as=1.44e-12 pd=6.96e-6 ps=6.96e-6 nrd=90e-3 nrs=90e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mnm5 net1 bias1 0 0 n18 m=1 w=w5 l=l5 nf=4 ad='w5/4<419.5e-9?(int(2.0)*(176.4e-15+(w5/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w5/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w5/4))+(2.0-int(2.0)!=0?480e-9*(w5/4):0))/1' as='w5/4<419.5e-9?((((176.4e-15+(w5/4)*100e-9)+0*(w5/4<419.5e-9?420e-9:w5/4))+int(1.5)*(176.4e-15+(w5/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w5/4)*100e-9:0))/1:(((480e-9*(w5/4)+0*(w5/4<419.5e-9?420e-9:w5/4))+int(1.5)*(540e-9*(w5/4)))+(2.0-int(2.0)==0?480e-9*(w5/4):0))/1' pd='w5/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w5/4))+(2.0-int(2.0)!=0?960e-9+2*(w5/4):0))/1' ps='w5/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w5/4))+0)+int(1.5)*(1.08e-6+2*(w5/4)))+(2.0-int(2.0)==0?960e-9+2*(w5/4):0))/1' nrd='270e-9/((w5/4)*4)' nrs='270e-9/((w5/4)*4)' sa='w5/4<419.5e-9?520e-9:480e-9' sb='w5/4<419.5e-9?520e-9:480e-9' sd='w5/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mnm4 vout net5 0 0 n18 m=1 w=w4 l=l4 nf=4 ad='w4/4<529.5e-9?(int(2.0)*(222.6e-15+(w4/4)*200e-9)+(2.0-int(2.0)!=0?222.6e-15+(w4/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w4/4))+(2.0-int(2.0)!=0?480e-9*(w4/4):0))/1' as='w4/4<529.5e-9?((((222.6e-15+(w4/4)*100e-9)+0*(w4/4<529.5e-9?530e-9:w4/4))+int(1.5)*(222.6e-15+(w4/4)*200e-9))+(2.0-int(2.0)==0?222.6e-15+(w4/4)*100e-9:0))/1:(((480e-9*(w4/4)+0*(w4/4<529.5e-9?530e-9:w4/4))+int(1.5)*(540e-9*(w4/4)))+(2.0-int(2.0)==0?480e-9*(w4/4):0))/1' pd='w4/4<529.5e-9?(int(2.0)*2.3e-6+(2.0-int(2.0)!=0?2.1e-6:0))/1:(int(2.0)*(1.08e-6+2*(w4/4))+(2.0-int(2.0)!=0?960e-9+2*(w4/4):0))/1' ps='w4/4<529.5e-9?((2.1e-6+int(1.5)*2.3e-6)+(2.0-int(2.0)==0?2.1e-6:0))/1:((((960e-9+2*(w4/4))+0)+int(1.5)*(1.08e-6+2*(w4/4)))+(2.0-int(2.0)==0?960e-9+2*(w4/4):0))/1' nrd='270e-9/((w4/4)*4)' nrs='270e-9/((w4/4)*4)' sa='w4/4<529.5e-9?520e-9:480e-9' sb='w4/4<529.5e-9?520e-9:480e-9' sd='w4/4<529.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mnm3 net5 net4 0 0 n18 m=1 w=w6 l=l6 nf=4 ad='w6/4<419.5e-9?(int(2.0)*(176.4e-15+(w6/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w6/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w6/4))+(2.0-int(2.0)!=0?480e-9*(w6/4):0))/1' as='w6/4<419.5e-9?((((176.4e-15+(w6/4)*100e-9)+0*(w6/4<419.5e-9?420e-9:w6/4))+int(1.5)*(176.4e-15+(w6/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w6/4)*100e-9:0))/1:(((480e-9*(w6/4)+0*(w6/4<419.5e-9?420e-9:w6/4))+int(1.5)*(540e-9*(w6/4)))+(2.0-int(2.0)==0?480e-9*(w6/4):0))/1' pd='w6/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w6/4))+(2.0-int(2.0)!=0?960e-9+2*(w6/4):0))/1' ps='w6/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w6/4))+0)+int(1.5)*(1.08e-6+2*(w6/4)))+(2.0-int(2.0)==0?960e-9+2*(w6/4):0))/1' nrd='270e-9/((w6/4)*4)' nrs='270e-9/((w6/4)*4)' sa='w6/4<419.5e-9?520e-9:480e-9' sb='w6/4<419.5e-9?520e-9:480e-9' sd='w6/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mnm2 net4 net4 0 0 n18 m=1 w=w6 l=l6 nf=4 ad='w6/4<529.5e-9?(int(2.0)*(222.6e-15+(w6/4)*200e-9)+(2.0-int(2.0)!=0?222.6e-15+(w6/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w6/4))+(2.0-int(2.0)!=0?480e-9*(w6/4):0))/1' as='w6/4<529.5e-9?((((222.6e-15+(w6/4)*100e-9)+0*(w6/4<529.5e-9?530e-9:w6/4))+int(1.5)*(222.6e-15+(w6/4)*200e-9))+(2.0-int(2.0)==0?222.6e-15+(w6/4)*100e-9:0))/1:(((480e-9*(w6/4)+0*(w6/4<529.5e-9?530e-9:w6/4))+int(1.5)*(540e-9*(w6/4)))+(2.0-int(2.0)==0?480e-9*(w6/4):0))/1' pd='w6/4<529.5e-9?(int(2.0)*2.3e-6+(2.0-int(2.0)!=0?2.1e-6:0))/1:(int(2.0)*(1.08e-6+2*(w6/4))+(2.0-int(2.0)!=0?960e-9+2*(w6/4):0))/1' ps='w6/4<529.5e-9?((2.1e-6+int(1.5)*2.3e-6)+(2.0-int(2.0)==0?2.1e-6:0))/1:((((960e-9+2*(w6/4))+0)+int(1.5)*(1.08e-6+2*(w6/4)))+(2.0-int(2.0)==0?960e-9+2*(w6/4):0))/1' nrd='270e-9/((w6/4)*4)' nrs='270e-9/((w6/4)*4)' sa='w6/4<529.5e-9?520e-9:480e-9' sb='w6/4<529.5e-9?520e-9:480e-9' sd='w6/4<529.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mnm1 net3 _net0 net1 0 n18 m=1 w=w2 l=l2 nf=4 ad='w2/4<419.5e-9?(int(2.0)*(176.4e-15+(w2/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w2/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w2/4))+(2.0-int(2.0)!=0?480e-9*(w2/4):0))/1' as='w2/4<419.5e-9?((((176.4e-15+(w2/4)*100e-9)+0*(w2/4<419.5e-9?420e-9:w2/4))+int(1.5)*(176.4e-15+(w2/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w2/4)*100e-9:0))/1:(((480e-9*(w2/4)+0*(w2/4<419.5e-9?420e-9:w2/4))+int(1.5)*(540e-9*(w2/4)))+(2.0-int(2.0)==0?480e-9*(w2/4):0))/1' pd='w2/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w2/4))+(2.0-int(2.0)!=0?960e-9+2*(w2/4):0))/1' ps='w2/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w2/4))+0)+int(1.5)*(1.08e-6+2*(w2/4)))+(2.0-int(2.0)==0?960e-9+2*(w2/4):0))/1' nrd='270e-9/((w2/4)*4)' nrs='270e-9/((w2/4)*4)' sa='w2/4<419.5e-9?520e-9:480e-9' sb='w2/4<419.5e-9?520e-9:480e-9' sd='w2/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mnm0 net2 _net1 net1 0 n18 m=1 w=w2 l=l2 nf=4 ad='w2/4<419.5e-9?(int(2.0)*(176.4e-15+(w2/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w2/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w2/4))+(2.0-int(2.0)!=0?480e-9*(w2/4):0))/1' as='w2/4<419.5e-9?((((176.4e-15+(w2/4)*100e-9)+0*(w2/4<419.5e-9?420e-9:w2/4))+int(1.5)*(176.4e-15+(w2/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w2/4)*100e-9:0))/1:(((480e-9*(w2/4)+0*(w2/4<419.5e-9?420e-9:w2/4))+int(1.5)*(540e-9*(w2/4)))+(2.0-int(2.0)==0?480e-9*(w2/4):0))/1' pd='w2/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w2/4))+(2.0-int(2.0)!=0?960e-9+2*(w2/4):0))/1' ps='w2/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w2/4))+0)+int(1.5)*(1.08e-6+2*(w2/4)))+(2.0-int(2.0)==0?960e-9+2*(w2/4):0))/1' nrd='270e-9/((w2/4)*4)' nrs='270e-9/((w2/4)*4)' sa='w2/4<419.5e-9?520e-9:480e-9' sb='w2/4<419.5e-9?520e-9:480e-9' sd='w2/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm7 bias3 bias3 vdd! vdd! p18 m=1 w=15e-6 l=1e-6 nf=1 ad=7.2e-12 as=7.2e-12 pd=30.96e-6 ps=30.96e-6 nrd=18e-3 nrs=18e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mpm5 bias2 bias2 vdd! vdd! p18 m=1 w=15e-6 l=1e-6 nf=1 ad=7.2e-12 as=7.2e-12 pd=30.96e-6 ps=30.96e-6 nrd=18e-3 nrs=18e-3 sa=480e-9 sb=480e-9 sd=0 sca=0 scb=0 scc=0
mpm4 vout bias3 vdd! vdd! p18 m=1 w=w8 l=l8 nf=4 ad='w8/4<419.5e-9?(int(2.0)*(176.4e-15+(w8/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w8/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w8/4))+(2.0-int(2.0)!=0?480e-9*(w8/4):0))/1' as='w8/4<419.5e-9?((((176.4e-15+(w8/4)*100e-9)+0*(w8/4<419.5e-9?420e-9:w8/4))+int(1.5)*(176.4e-15+(w8/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w8/4)*100e-9:0))/1:(((480e-9*(w8/4)+0*(w8/4<419.5e-9?420e-9:w8/4))+int(1.5)*(540e-9*(w8/4)))+(2.0-int(2.0)==0?480e-9*(w8/4):0))/1' pd='w8/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w8/4))+(2.0-int(2.0)!=0?960e-9+2*(w8/4):0))/1' ps='w8/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w8/4))+0)+int(1.5)*(1.08e-6+2*(w8/4)))+(2.0-int(2.0)==0?960e-9+2*(w8/4):0))/1' nrd='270e-9/((w8/4)*4)' nrs='270e-9/((w8/4)*4)' sa='w8/4<419.5e-9?520e-9:480e-9' sb='w8/4<419.5e-9?520e-9:480e-9' sd='w8/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm3 net5 bias2 vdd! vdd! p18 m=1 w=w7 l=l7 nf=4 ad='w7/4<419.5e-9?(int(2.0)*(176.4e-15+(w7/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w7/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w7/4))+(2.0-int(2.0)!=0?480e-9*(w7/4):0))/1' as='w7/4<419.5e-9?((((176.4e-15+(w7/4)*100e-9)+0*(w7/4<419.5e-9?420e-9:w7/4))+int(1.5)*(176.4e-15+(w7/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w7/4)*100e-9:0))/1:(((480e-9*(w7/4)+0*(w7/4<419.5e-9?420e-9:w7/4))+int(1.5)*(540e-9*(w7/4)))+(2.0-int(2.0)==0?480e-9*(w7/4):0))/1' pd='w7/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w7/4))+(2.0-int(2.0)!=0?960e-9+2*(w7/4):0))/1' ps='w7/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w7/4))+0)+int(1.5)*(1.08e-6+2*(w7/4)))+(2.0-int(2.0)==0?960e-9+2*(w7/4):0))/1' nrd='270e-9/((w7/4)*4)' nrs='270e-9/((w7/4)*4)' sa='w7/4<419.5e-9?520e-9:480e-9' sb='w7/4<419.5e-9?520e-9:480e-9' sd='w7/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm2 net4 net3 vdd! vdd! p18 m=1 w=w3 l=l3 nf=4 ad='w3/4<419.5e-9?(int(2.0)*(176.4e-15+(w3/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w3/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w3/4))+(2.0-int(2.0)!=0?480e-9*(w3/4):0))/1' as='w3/4<419.5e-9?((((176.4e-15+(w3/4)*100e-9)+0*(w3/4<419.5e-9?420e-9:w3/4))+int(1.5)*(176.4e-15+(w3/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w3/4)*100e-9:0))/1:(((480e-9*(w3/4)+0*(w3/4<419.5e-9?420e-9:w3/4))+int(1.5)*(540e-9*(w3/4)))+(2.0-int(2.0)==0?480e-9*(w3/4):0))/1' pd='w3/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w3/4))+(2.0-int(2.0)!=0?960e-9+2*(w3/4):0))/1' ps='w3/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w3/4))+0)+int(1.5)*(1.08e-6+2*(w3/4)))+(2.0-int(2.0)==0?960e-9+2*(w3/4):0))/1' nrd='270e-9/((w3/4)*4)' nrs='270e-9/((w3/4)*4)' sa='w3/4<419.5e-9?520e-9:480e-9' sb='w3/4<419.5e-9?520e-9:480e-9' sd='w3/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm1 net2 net2 vdd! vdd! p18 m=1 w=w1 l=l1 nf=4 ad='w1/4<419.5e-9?(int(2.0)*(176.4e-15+(w1/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w1/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w1/4))+(2.0-int(2.0)!=0?480e-9*(w1/4):0))/1' as='w1/4<419.5e-9?((((176.4e-15+(w1/4)*100e-9)+0*(w1/4<419.5e-9?420e-9:w1/4))+int(1.5)*(176.4e-15+(w1/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w1/4)*100e-9:0))/1:(((480e-9*(w1/4)+0*(w1/4<419.5e-9?420e-9:w1/4))+int(1.5)*(540e-9*(w1/4)))+(2.0-int(2.0)==0?480e-9*(w1/4):0))/1' pd='w1/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w1/4))+(2.0-int(2.0)!=0?960e-9+2*(w1/4):0))/1' ps='w1/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w1/4))+0)+int(1.5)*(1.08e-6+2*(w1/4)))+(2.0-int(2.0)==0?960e-9+2*(w1/4):0))/1' nrd='270e-9/((w1/4)*4)' nrs='270e-9/((w1/4)*4)' sa='w1/4<419.5e-9?520e-9:480e-9' sb='w1/4<419.5e-9?520e-9:480e-9' sd='w1/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
mpm0 net3 net2 vdd! vdd! p18 m=1 w=w1 l=l1 nf=4 ad='w1/4<419.5e-9?(int(2.0)*(176.4e-15+(w1/4)*200e-9)+(2.0-int(2.0)!=0?176.4e-15+(w1/4)*100e-9:0))/1:(int(2.0)*(540e-9*(w1/4))+(2.0-int(2.0)!=0?480e-9*(w1/4):0))/1' as='w1/4<419.5e-9?((((176.4e-15+(w1/4)*100e-9)+0*(w1/4<419.5e-9?420e-9:w1/4))+int(1.5)*(176.4e-15+(w1/4)*200e-9))+(2.0-int(2.0)==0?176.4e-15+(w1/4)*100e-9:0))/1:(((480e-9*(w1/4)+0*(w1/4<419.5e-9?420e-9:w1/4))+int(1.5)*(540e-9*(w1/4)))+(2.0-int(2.0)==0?480e-9*(w1/4):0))/1' pd='w1/4<419.5e-9?(int(2.0)*2.08e-6+(2.0-int(2.0)!=0?1.88e-6:0))/1:(int(2.0)*(1.08e-6+2*(w1/4))+(2.0-int(2.0)!=0?960e-9+2*(w1/4):0))/1' ps='w1/4<419.5e-9?((1.88e-6+int(1.5)*2.08e-6)+(2.0-int(2.0)==0?1.88e-6:0))/1:((((960e-9+2*(w1/4))+0)+int(1.5)*(1.08e-6+2*(w1/4)))+(2.0-int(2.0)==0?960e-9+2*(w1/4):0))/1' nrd='270e-9/((w1/4)*4)' nrs='270e-9/((w1/4)*4)' sa='w1/4<419.5e-9?520e-9:480e-9' sb='w1/4<419.5e-9?520e-9:480e-9' sd='w1/4<419.5e-9?620e-9:540e-9' sca=0 scb=0 scc=0
c1 net3 vout c1
c0 net5 vout c2
i6 bias3 0 DC=20e-6
i3 bias2 0 DC=20e-6
i2 vdd! bias1 DC=20e-6
.ends OTA_three
** End of subcircuit definition.

** Library name: ZYX_try
** Cell name: tb_OTA_three
** View name: schematic
xi0 net2 net3 net1 OTA_three
v9 net3 0 DC=900e-3 AC 0 0
v2 vdd! 0 DC=1.8
v6 net2 net1 DC=0 AC 1 180
c0 net1 0 5e-12

.control
op
AC DEC 10 0.01 100000K
.endc

.END
